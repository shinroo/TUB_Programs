library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bin2Char is
	port(bin : in std_logic_vector(3 downto 0);
		 bitmask : out std_logic_vector(6 downto 0));
end bin2Char;

architecture behavioral of bin2Char is   
begin
	
	-- bin2Char-Beschreibung hier einfügen
	 
end behavioral;
