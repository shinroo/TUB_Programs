library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity reg is
	generic(
		WIDTH : integer);
	port(
		clk : in  std_logic;
		rst : in  std_logic;
		en  : in  std_logic;
		D   : in  std_logic_vector( WIDTH - 1 downto 0 );
		Q   : out std_logic_vector( WIDTH - 1 downto 0 ));
end reg;

architecture behavioral of reg is
begin
	process (clk)
	variable i : integer := WIDTH - 1;
	variable temp : std_logic_vector(WIDTH - 1 downto 0) := (others => '0');
	begin
		if (clk = '1' and clk'last_value = '0' and rst = '1') then
			Q <= (others => '0');
		elsif (clk = '1' and clk'last_value = '0' and en = '1') then
			Q <= D;
		end if;
	end process;
	
end behavioral;
